`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:02:15 10/10/2015 
// Design Name: 
// Module Name:    neg2pos 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module neg2pos(
    input [15:0] i,
    output [15:0] o
    );
	 
	 reg[15:0] interm;
	 
	 // Signed Adder
	 
	 always@(*) begin
		
	 end
	 
endmodule
